package words_lengths_pkg;

    parameter integer Nsig = 3; //Number bits of signal
    parameter integer Ncoef = 3; //Number bits of coefficients
    parameter integer Nstage = 3; //Number of stages

endpackage
